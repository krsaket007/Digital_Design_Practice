VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO MUX_2X1
   CLASS BLOCK ;
   FOREIGN MUX_2X1 ;
   ORIGIN 2.6000 -0.0000 ;
   SIZE 18.7000 BY 11.0000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.6000 0.8000 1.0000 3.1000 ;
	    RECT 3.8000 0.8000 4.2000 5.1000 ;
	    RECT 5.9000 0.8000 6.3000 3.1000 ;
	    RECT 7.0000 0.8000 7.4000 3.1000 ;
	    RECT 8.6000 0.8000 9.0000 3.1000 ;
	    RECT 11.8000 0.8000 12.2000 4.5000 ;
	    RECT 0.2000 0.2000 13.4000 0.8000 ;
         LAYER metal2 ;
	    RECT 1.6000 0.3000 3.2000 0.7000 ;
         LAYER metal3 ;
	    RECT 1.6000 0.3000 3.2000 0.7000 ;
         LAYER metal4 ;
	    RECT 1.6000 0.3000 3.2000 0.7000 ;
         LAYER metal5 ;
	    RECT 1.6000 0.7000 2.2000 0.8000 ;
	    RECT 2.6000 0.7000 3.2000 0.8000 ;
	    RECT 1.6000 0.2000 3.2000 0.7000 ;
         LAYER metal6 ;
	    RECT 1.6000 0.0000 3.2000 11.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 10.2000 13.4000 10.8000 ;
	    RECT 0.6000 8.9000 1.0000 10.2000 ;
	    RECT 4.6000 8.3000 5.0000 10.2000 ;
	    RECT 8.6000 7.9000 9.0000 10.2000 ;
	    RECT 11.8000 7.9000 12.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 8.8000 10.3000 10.4000 10.7000 ;
         LAYER metal3 ;
	    RECT 8.8000 10.3000 10.4000 10.7000 ;
         LAYER metal4 ;
	    RECT 8.8000 10.3000 10.4000 10.7000 ;
         LAYER metal5 ;
	    RECT 8.8000 10.7000 9.4000 10.8000 ;
	    RECT 9.8000 10.7000 10.4000 10.8000 ;
	    RECT 8.8000 10.2000 10.4000 10.7000 ;
         LAYER metal6 ;
	    RECT 8.8000 0.0000 10.4000 11.0000 ;
      END
   END gnd
   PIN inp_1
      PORT
         LAYER metal1 ;
	    RECT 0.6000 7.8000 1.0000 8.6000 ;
	    RECT 0.6000 7.2000 0.9000 7.8000 ;
	    RECT 0.6000 6.8000 1.0000 7.2000 ;
         LAYER metal2 ;
	    RECT 0.6000 7.8000 1.0000 8.2000 ;
	    RECT 0.6000 7.2000 0.9000 7.8000 ;
	    RECT 0.6000 6.8000 1.0000 7.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 8.1000 1.0000 8.2000 ;
	    RECT -2.6000 7.8000 1.0000 8.1000 ;
      END
   END inp_1
   PIN inp_2
      PORT
         LAYER metal1 ;
	    RECT 8.6000 7.1000 9.0000 7.6000 ;
	    RECT 10.2000 7.1000 10.6000 7.2000 ;
	    RECT 8.6000 6.8000 10.6000 7.1000 ;
         LAYER metal2 ;
	    RECT 10.2000 7.8000 10.6000 8.2000 ;
	    RECT 10.2000 7.2000 10.5000 7.8000 ;
	    RECT 10.2000 6.8000 10.6000 7.2000 ;
         LAYER metal3 ;
	    RECT 10.2000 8.1000 10.6000 8.2000 ;
	    RECT 10.2000 7.8000 16.1000 8.1000 ;
      END
   END inp_2
   PIN sel
      PORT
         LAYER metal1 ;
	    RECT 4.6000 5.8000 5.0000 6.6000 ;
	    RECT 7.0000 4.4000 7.4000 5.2000 ;
         LAYER metal2 ;
	    RECT 4.6000 6.8000 5.0000 7.2000 ;
	    RECT 4.6000 6.2000 4.9000 6.8000 ;
	    RECT 4.6000 5.8000 5.0000 6.2000 ;
	    RECT 7.0000 5.8000 7.4000 6.2000 ;
	    RECT 7.0000 5.2000 7.3000 5.8000 ;
	    RECT 7.0000 4.8000 7.4000 5.2000 ;
         LAYER metal3 ;
	    RECT 4.6000 6.8000 5.0000 7.2000 ;
	    RECT 4.6000 6.1000 4.9000 6.8000 ;
	    RECT 7.0000 6.1000 7.4000 6.2000 ;
	    RECT -2.6000 5.8000 7.4000 6.1000 ;
      END
   END sel
   PIN out
      PORT
         LAYER metal1 ;
	    RECT 12.6000 6.2000 13.0000 9.9000 ;
	    RECT 12.7000 5.1000 13.0000 6.2000 ;
	    RECT 12.6000 1.1000 13.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 12.6000 6.8000 13.0000 7.2000 ;
	    RECT 12.6000 6.2000 12.9000 6.8000 ;
	    RECT 12.6000 5.8000 13.0000 6.2000 ;
         LAYER metal3 ;
	    RECT 12.6000 6.1000 13.0000 6.2000 ;
	    RECT 12.6000 5.8000 16.1000 6.1000 ;
      END
   END out
   OBS
         LAYER metal1 ;
	    RECT 1.4000 7.1000 1.8000 9.9000 ;
	    RECT 3.8000 8.0000 4.2000 9.9000 ;
	    RECT 5.4000 8.0000 5.8000 9.9000 ;
	    RECT 3.8000 7.9000 5.8000 8.0000 ;
	    RECT 6.2000 7.9000 6.6000 9.9000 ;
	    RECT 7.3000 8.2000 7.7000 9.9000 ;
	    RECT 7.3000 7.9000 8.2000 8.2000 ;
	    RECT 3.9000 7.7000 5.7000 7.9000 ;
	    RECT 4.2000 7.2000 4.6000 7.4000 ;
	    RECT 6.2000 7.2000 6.5000 7.9000 ;
	    RECT 3.8000 7.1000 4.6000 7.2000 ;
	    RECT 1.4000 6.9000 4.6000 7.1000 ;
	    RECT 5.3000 7.1000 6.6000 7.2000 ;
	    RECT 7.0000 7.1000 7.4000 7.2000 ;
	    RECT 1.4000 6.8000 4.2000 6.9000 ;
	    RECT 5.3000 6.8000 7.4000 7.1000 ;
	    RECT 1.4000 1.1000 1.8000 6.8000 ;
	    RECT 5.3000 5.1000 5.6000 6.8000 ;
	    RECT 7.8000 6.1000 8.2000 7.9000 ;
	    RECT 11.0000 7.6000 11.4000 9.9000 ;
	    RECT 11.0000 7.3000 12.1000 7.6000 ;
	    RECT 6.2000 5.8000 8.2000 6.1000 ;
	    RECT 11.0000 5.8000 11.4000 6.6000 ;
	    RECT 11.8000 5.8000 12.1000 7.3000 ;
	    RECT 6.2000 5.2000 6.5000 5.8000 ;
	    RECT 6.2000 5.1000 6.6000 5.2000 ;
	    RECT 5.1000 4.8000 5.6000 5.1000 ;
	    RECT 5.9000 4.8000 6.6000 5.1000 ;
	    RECT 5.1000 1.1000 5.5000 4.8000 ;
	    RECT 5.9000 4.2000 6.2000 4.8000 ;
	    RECT 5.8000 3.8000 6.2000 4.2000 ;
	    RECT 7.8000 1.1000 8.2000 5.8000 ;
	    RECT 11.8000 5.4000 12.4000 5.8000 ;
	    RECT 11.8000 5.1000 12.1000 5.4000 ;
	    RECT 11.0000 4.8000 12.1000 5.1000 ;
	    RECT 11.0000 1.1000 11.4000 4.8000 ;
         LAYER metal2 ;
	    RECT 6.2000 7.1000 6.6000 7.2000 ;
	    RECT 7.0000 7.1000 7.4000 7.2000 ;
	    RECT 6.2000 6.8000 7.4000 7.1000 ;
	    RECT 11.0000 6.8000 11.4000 7.2000 ;
	    RECT 11.0000 6.2000 11.3000 6.8000 ;
	    RECT 11.0000 5.8000 11.4000 6.2000 ;
         LAYER metal3 ;
	    RECT 6.2000 7.1000 6.6000 7.2000 ;
	    RECT 11.0000 7.1000 11.4000 7.2000 ;
	    RECT 6.2000 6.8000 11.4000 7.1000 ;
   END
END MUX_2X1
